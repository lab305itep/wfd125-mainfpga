localparam VERSION = 32'h00020003;