localparam VERSION = 32'h00020001;